module matdet10 #(parameter DATA_WIDTH=8, parameter MATRIX_SIZE=100) (input wire [(MATRIX_SIZE * DATA_WIDTH) - 1:0] a, output wire [DATA_WIDTH-1:0] det);
wire [DATA_WIDTH-1:0] w0, w1, w2, w3, w4, w5, w6, w7, w8, w9, w10, w11, w12, w13, w14, w15, w16, w17, w18, w19, w20, w21, w22, w23, w24, w25, w26, w27, w28;
matdet9 md0({a[95:88], a[103:96], a[111:104], a[119:112], a[127:120], a[135:128], a[143:136], a[151:144], a[159:152], a[175:168], a[183:176], a[191:184], a[199:192], a[207:200], a[215:208], a[223:216], a[231:224], a[239:232], a[255:248], a[263:256], a[271:264], a[279:272], a[287:280], a[295:288], a[303:296], a[311:304], a[319:312], a[335:328], a[343:336], a[351:344], a[359:352], a[367:360], a[375:368], a[383:376], a[391:384], a[399:392], a[415:408], a[423:416], a[431:424], a[439:432], a[447:440], a[455:448], a[463:456], a[471:464], a[479:472], a[495:488], a[503:496], a[511:504], a[519:512], a[527:520], a[535:528], a[543:536], a[551:544], a[559:552], a[575:568], a[583:576], a[591:584], a[599:592], a[607:600], a[615:608], a[623:616], a[631:624], a[639:632], a[655:648], a[663:656], a[671:664], a[679:672], a[687:680], a[695:688], a[703:696], a[711:704], a[719:712], a[735:728], a[743:736], a[751:744], a[759:752], a[767:760], a[775:768], a[783:776], a[791:784], a[799:792]}, w0);
matdet9 md1({a[87:80], a[103:96], a[111:104], a[119:112], a[127:120], a[135:128], a[143:136], a[151:144], a[159:152], a[167:160], a[183:176], a[191:184], a[199:192], a[207:200], a[215:208], a[223:216], a[231:224], a[239:232], a[247:240], a[263:256], a[271:264], a[279:272], a[287:280], a[295:288], a[303:296], a[311:304], a[319:312], a[327:320], a[343:336], a[351:344], a[359:352], a[367:360], a[375:368], a[383:376], a[391:384], a[399:392], a[407:400], a[423:416], a[431:424], a[439:432], a[447:440], a[455:448], a[463:456], a[471:464], a[479:472], a[487:480], a[503:496], a[511:504], a[519:512], a[527:520], a[535:528], a[543:536], a[551:544], a[559:552], a[567:560], a[583:576], a[591:584], a[599:592], a[607:600], a[615:608], a[623:616], a[631:624], a[639:632], a[647:640], a[663:656], a[671:664], a[679:672], a[687:680], a[695:688], a[703:696], a[711:704], a[719:712], a[727:720], a[743:736], a[751:744], a[759:752], a[767:760], a[775:768], a[783:776], a[791:784], a[799:792]}, w1);
matdet9 md2({a[87:80], a[95:88], a[111:104], a[119:112], a[127:120], a[135:128], a[143:136], a[151:144], a[159:152], a[167:160], a[175:168], a[191:184], a[199:192], a[207:200], a[215:208], a[223:216], a[231:224], a[239:232], a[247:240], a[255:248], a[271:264], a[279:272], a[287:280], a[295:288], a[303:296], a[311:304], a[319:312], a[327:320], a[335:328], a[351:344], a[359:352], a[367:360], a[375:368], a[383:376], a[391:384], a[399:392], a[407:400], a[415:408], a[431:424], a[439:432], a[447:440], a[455:448], a[463:456], a[471:464], a[479:472], a[487:480], a[495:488], a[511:504], a[519:512], a[527:520], a[535:528], a[543:536], a[551:544], a[559:552], a[567:560], a[575:568], a[591:584], a[599:592], a[607:600], a[615:608], a[623:616], a[631:624], a[639:632], a[647:640], a[655:648], a[671:664], a[679:672], a[687:680], a[695:688], a[703:696], a[711:704], a[719:712], a[727:720], a[735:728], a[751:744], a[759:752], a[767:760], a[775:768], a[783:776], a[791:784], a[799:792]}, w2);
matdet9 md3({a[87:80], a[95:88], a[103:96], a[119:112], a[127:120], a[135:128], a[143:136], a[151:144], a[159:152], a[167:160], a[175:168], a[183:176], a[199:192], a[207:200], a[215:208], a[223:216], a[231:224], a[239:232], a[247:240], a[255:248], a[263:256], a[279:272], a[287:280], a[295:288], a[303:296], a[311:304], a[319:312], a[327:320], a[335:328], a[343:336], a[359:352], a[367:360], a[375:368], a[383:376], a[391:384], a[399:392], a[407:400], a[415:408], a[423:416], a[439:432], a[447:440], a[455:448], a[463:456], a[471:464], a[479:472], a[487:480], a[495:488], a[503:496], a[519:512], a[527:520], a[535:528], a[543:536], a[551:544], a[559:552], a[567:560], a[575:568], a[583:576], a[599:592], a[607:600], a[615:608], a[623:616], a[631:624], a[639:632], a[647:640], a[655:648], a[663:656], a[679:672], a[687:680], a[695:688], a[703:696], a[711:704], a[719:712], a[727:720], a[735:728], a[743:736], a[759:752], a[767:760], a[775:768], a[783:776], a[791:784], a[799:792]}, w3);
matdet9 md4({a[87:80], a[95:88], a[103:96], a[111:104], a[127:120], a[135:128], a[143:136], a[151:144], a[159:152], a[167:160], a[175:168], a[183:176], a[191:184], a[207:200], a[215:208], a[223:216], a[231:224], a[239:232], a[247:240], a[255:248], a[263:256], a[271:264], a[287:280], a[295:288], a[303:296], a[311:304], a[319:312], a[327:320], a[335:328], a[343:336], a[351:344], a[367:360], a[375:368], a[383:376], a[391:384], a[399:392], a[407:400], a[415:408], a[423:416], a[431:424], a[447:440], a[455:448], a[463:456], a[471:464], a[479:472], a[487:480], a[495:488], a[503:496], a[511:504], a[527:520], a[535:528], a[543:536], a[551:544], a[559:552], a[567:560], a[575:568], a[583:576], a[591:584], a[607:600], a[615:608], a[623:616], a[631:624], a[639:632], a[647:640], a[655:648], a[663:656], a[671:664], a[687:680], a[695:688], a[703:696], a[711:704], a[719:712], a[727:720], a[735:728], a[743:736], a[751:744], a[767:760], a[775:768], a[783:776], a[791:784], a[799:792]}, w4);
matdet9 md5({a[87:80], a[95:88], a[103:96], a[111:104], a[119:112], a[135:128], a[143:136], a[151:144], a[159:152], a[167:160], a[175:168], a[183:176], a[191:184], a[199:192], a[215:208], a[223:216], a[231:224], a[239:232], a[247:240], a[255:248], a[263:256], a[271:264], a[279:272], a[295:288], a[303:296], a[311:304], a[319:312], a[327:320], a[335:328], a[343:336], a[351:344], a[359:352], a[375:368], a[383:376], a[391:384], a[399:392], a[407:400], a[415:408], a[423:416], a[431:424], a[439:432], a[455:448], a[463:456], a[471:464], a[479:472], a[487:480], a[495:488], a[503:496], a[511:504], a[519:512], a[535:528], a[543:536], a[551:544], a[559:552], a[567:560], a[575:568], a[583:576], a[591:584], a[599:592], a[615:608], a[623:616], a[631:624], a[639:632], a[647:640], a[655:648], a[663:656], a[671:664], a[679:672], a[695:688], a[703:696], a[711:704], a[719:712], a[727:720], a[735:728], a[743:736], a[751:744], a[759:752], a[775:768], a[783:776], a[791:784], a[799:792]}, w5);
matdet9 md6({a[87:80], a[95:88], a[103:96], a[111:104], a[119:112], a[127:120], a[143:136], a[151:144], a[159:152], a[167:160], a[175:168], a[183:176], a[191:184], a[199:192], a[207:200], a[223:216], a[231:224], a[239:232], a[247:240], a[255:248], a[263:256], a[271:264], a[279:272], a[287:280], a[303:296], a[311:304], a[319:312], a[327:320], a[335:328], a[343:336], a[351:344], a[359:352], a[367:360], a[383:376], a[391:384], a[399:392], a[407:400], a[415:408], a[423:416], a[431:424], a[439:432], a[447:440], a[463:456], a[471:464], a[479:472], a[487:480], a[495:488], a[503:496], a[511:504], a[519:512], a[527:520], a[543:536], a[551:544], a[559:552], a[567:560], a[575:568], a[583:576], a[591:584], a[599:592], a[607:600], a[623:616], a[631:624], a[639:632], a[647:640], a[655:648], a[663:656], a[671:664], a[679:672], a[687:680], a[703:696], a[711:704], a[719:712], a[727:720], a[735:728], a[743:736], a[751:744], a[759:752], a[767:760], a[783:776], a[791:784], a[799:792]}, w6);
matdet9 md7({a[87:80], a[95:88], a[103:96], a[111:104], a[119:112], a[127:120], a[135:128], a[151:144], a[159:152], a[167:160], a[175:168], a[183:176], a[191:184], a[199:192], a[207:200], a[215:208], a[231:224], a[239:232], a[247:240], a[255:248], a[263:256], a[271:264], a[279:272], a[287:280], a[295:288], a[311:304], a[319:312], a[327:320], a[335:328], a[343:336], a[351:344], a[359:352], a[367:360], a[375:368], a[391:384], a[399:392], a[407:400], a[415:408], a[423:416], a[431:424], a[439:432], a[447:440], a[455:448], a[471:464], a[479:472], a[487:480], a[495:488], a[503:496], a[511:504], a[519:512], a[527:520], a[535:528], a[551:544], a[559:552], a[567:560], a[575:568], a[583:576], a[591:584], a[599:592], a[607:600], a[615:608], a[631:624], a[639:632], a[647:640], a[655:648], a[663:656], a[671:664], a[679:672], a[687:680], a[695:688], a[711:704], a[719:712], a[727:720], a[735:728], a[743:736], a[751:744], a[759:752], a[767:760], a[775:768], a[791:784], a[799:792]}, w7);
matdet9 md8({a[87:80], a[95:88], a[103:96], a[111:104], a[119:112], a[127:120], a[135:128], a[143:136], a[159:152], a[167:160], a[175:168], a[183:176], a[191:184], a[199:192], a[207:200], a[215:208], a[223:216], a[239:232], a[247:240], a[255:248], a[263:256], a[271:264], a[279:272], a[287:280], a[295:288], a[303:296], a[319:312], a[327:320], a[335:328], a[343:336], a[351:344], a[359:352], a[367:360], a[375:368], a[383:376], a[399:392], a[407:400], a[415:408], a[423:416], a[431:424], a[439:432], a[447:440], a[455:448], a[463:456], a[479:472], a[487:480], a[495:488], a[503:496], a[511:504], a[519:512], a[527:520], a[535:528], a[543:536], a[559:552], a[567:560], a[575:568], a[583:576], a[591:584], a[599:592], a[607:600], a[615:608], a[623:616], a[639:632], a[647:640], a[655:648], a[663:656], a[671:664], a[679:672], a[687:680], a[695:688], a[703:696], a[719:712], a[727:720], a[735:728], a[743:736], a[751:744], a[759:752], a[767:760], a[775:768], a[783:776], a[799:792]}, w8);
matdet9 md9({a[87:80], a[95:88], a[103:96], a[111:104], a[119:112], a[127:120], a[135:128], a[143:136], a[151:144], a[167:160], a[175:168], a[183:176], a[191:184], a[199:192], a[207:200], a[215:208], a[223:216], a[231:224], a[247:240], a[255:248], a[263:256], a[271:264], a[279:272], a[287:280], a[295:288], a[303:296], a[311:304], a[327:320], a[335:328], a[343:336], a[351:344], a[359:352], a[367:360], a[375:368], a[383:376], a[391:384], a[407:400], a[415:408], a[423:416], a[431:424], a[439:432], a[447:440], a[455:448], a[463:456], a[471:464], a[487:480], a[495:488], a[503:496], a[511:504], a[519:512], a[527:520], a[535:528], a[543:536], a[551:544], a[567:560], a[575:568], a[583:576], a[591:584], a[599:592], a[607:600], a[615:608], a[623:616], a[631:624], a[647:640], a[655:648], a[663:656], a[671:664], a[679:672], a[687:680], a[695:688], a[703:696], a[711:704], a[727:720], a[735:728], a[743:736], a[751:744], a[759:752], a[767:760], a[775:768], a[783:776], a[791:784]}, w9);
mul m0(a[7:0], w0, w10);
mul m1(a[15:8], w1, w11);
mul m2(a[23:16], w2, w12);
mul m3(a[31:24], w3, w13);
mul m4(a[39:32], w4, w14);
mul m5(a[47:40], w5, w15);
mul m6(a[55:48], w6, w16);
mul m7(a[63:56], w7, w17);
mul m8(a[71:64], w8, w18);
mul m9(a[79:72], w9, w19);
sub op0(w10, w11, w20);
add op1(w20, w12, w21);
sub op2(w21, w13, w22);
add op3(w22, w14, w23);
sub op4(w23, w15, w24);
add op5(w24, w16, w25);
sub op6(w25, w17, w26);
add op7(w26, w18, w27);
sub op8(w27, w19, det);
endmodule
