module matdet6 #(parameter DATA_WIDTH=8, parameter MATRIX_SIZE=36) (input wire [(MATRIX_SIZE * DATA_WIDTH) - 1:0] a, output wire [DATA_WIDTH-1:0] det);
wire [DATA_WIDTH-1:0] w0, w1, w2, w3, w4, w5, w6, w7, w8, w9, w10, w11, w12, w13, w14, w15, w16;
matdet5 md0({a[63:56], a[71:64], a[79:72], a[87:80], a[95:88], a[111:104], a[119:112], a[127:120], a[135:128], a[143:136], a[159:152], a[167:160], a[175:168], a[183:176], a[191:184], a[207:200], a[215:208], a[223:216], a[231:224], a[239:232], a[255:248], a[263:256], a[271:264], a[279:272], a[287:280]}, w0);
matdet5 md1({a[55:48], a[71:64], a[79:72], a[87:80], a[95:88], a[103:96], a[119:112], a[127:120], a[135:128], a[143:136], a[151:144], a[167:160], a[175:168], a[183:176], a[191:184], a[199:192], a[215:208], a[223:216], a[231:224], a[239:232], a[247:240], a[263:256], a[271:264], a[279:272], a[287:280]}, w1);
matdet5 md2({a[55:48], a[63:56], a[79:72], a[87:80], a[95:88], a[103:96], a[111:104], a[127:120], a[135:128], a[143:136], a[151:144], a[159:152], a[175:168], a[183:176], a[191:184], a[199:192], a[207:200], a[223:216], a[231:224], a[239:232], a[247:240], a[255:248], a[271:264], a[279:272], a[287:280]}, w2);
matdet5 md3({a[55:48], a[63:56], a[71:64], a[87:80], a[95:88], a[103:96], a[111:104], a[119:112], a[135:128], a[143:136], a[151:144], a[159:152], a[167:160], a[183:176], a[191:184], a[199:192], a[207:200], a[215:208], a[231:224], a[239:232], a[247:240], a[255:248], a[263:256], a[279:272], a[287:280]}, w3);
matdet5 md4({a[55:48], a[63:56], a[71:64], a[79:72], a[95:88], a[103:96], a[111:104], a[119:112], a[127:120], a[143:136], a[151:144], a[159:152], a[167:160], a[175:168], a[191:184], a[199:192], a[207:200], a[215:208], a[223:216], a[239:232], a[247:240], a[255:248], a[263:256], a[271:264], a[287:280]}, w4);
matdet5 md5({a[55:48], a[63:56], a[71:64], a[79:72], a[87:80], a[103:96], a[111:104], a[119:112], a[127:120], a[135:128], a[151:144], a[159:152], a[167:160], a[175:168], a[183:176], a[199:192], a[207:200], a[215:208], a[223:216], a[231:224], a[247:240], a[255:248], a[263:256], a[271:264], a[279:272]}, w5);
mul m0(a[7:0], w0, w6);
mul m1(a[15:8], w1, w7);
mul m2(a[23:16], w2, w8);
mul m3(a[31:24], w3, w9);
mul m4(a[39:32], w4, w10);
mul m5(a[47:40], w5, w11);
sub op0(w6, w7, w12);
add op1(w12, w8, w13);
sub op2(w13, w9, w14);
add op3(w14, w10, w15);
sub op4(w15, w11, det);
endmodule
