module matdet5 #(parameter DATA_WIDTH=8, parameter MATRIX_SIZE=25) (input wire [(MATRIX_SIZE * DATA_WIDTH) - 1:0] a, output wire [DATA_WIDTH-1:0] det);
wire [DATA_WIDTH-1:0] w0, w1, w2, w3, w4, w5, w6, w7, w8, w9, w10, w11, w12, w13;
matdet4 md0({a[55:48], a[63:56], a[71:64], a[79:72], a[95:88], a[103:96], a[111:104], a[119:112], a[135:128], a[143:136], a[151:144], a[159:152], a[175:168], a[183:176], a[191:184], a[199:192]}, w0);
matdet4 md1({a[47:40], a[63:56], a[71:64], a[79:72], a[87:80], a[103:96], a[111:104], a[119:112], a[127:120], a[143:136], a[151:144], a[159:152], a[167:160], a[183:176], a[191:184], a[199:192]}, w1);
matdet4 md2({a[47:40], a[55:48], a[71:64], a[79:72], a[87:80], a[95:88], a[111:104], a[119:112], a[127:120], a[135:128], a[151:144], a[159:152], a[167:160], a[175:168], a[191:184], a[199:192]}, w2);
matdet4 md3({a[47:40], a[55:48], a[63:56], a[79:72], a[87:80], a[95:88], a[103:96], a[119:112], a[127:120], a[135:128], a[143:136], a[159:152], a[167:160], a[175:168], a[183:176], a[199:192]}, w3);
matdet4 md4({a[47:40], a[55:48], a[63:56], a[71:64], a[87:80], a[95:88], a[103:96], a[111:104], a[127:120], a[135:128], a[143:136], a[151:144], a[167:160], a[175:168], a[183:176], a[191:184]}, w4);
mul m0(a[7:0], w0, w5);
mul m1(a[15:8], w1, w6);
mul m2(a[23:16], w2, w7);
mul m3(a[31:24], w3, w8);
mul m4(a[39:32], w4, w9);
sub op0(w5, w6, w10);
add op1(w10, w7, w11);
sub op2(w11, w8, w12);
add op3(w12, w9, det);
endmodule
