module matdet7 #(parameter DATA_WIDTH=8, parameter MATRIX_SIZE=49) (input wire [(MATRIX_SIZE * DATA_WIDTH) - 1:0] a, output wire [DATA_WIDTH-1:0] det);
wire [DATA_WIDTH-1:0] w0, w1, w2, w3, w4, w5, w6, w7, w8, w9, w10, w11, w12, w13, w14, w15, w16, w17, w18, w19;
matdet6 md0({a[71:64], a[79:72], a[87:80], a[95:88], a[103:96], a[111:104], a[127:120], a[135:128], a[143:136], a[151:144], a[159:152], a[167:160], a[183:176], a[191:184], a[199:192], a[207:200], a[215:208], a[223:216], a[239:232], a[247:240], a[255:248], a[263:256], a[271:264], a[279:272], a[295:288], a[303:296], a[311:304], a[319:312], a[327:320], a[335:328], a[351:344], a[359:352], a[367:360], a[375:368], a[383:376], a[391:384]}, w0);
matdet6 md1({a[63:56], a[79:72], a[87:80], a[95:88], a[103:96], a[111:104], a[119:112], a[135:128], a[143:136], a[151:144], a[159:152], a[167:160], a[175:168], a[191:184], a[199:192], a[207:200], a[215:208], a[223:216], a[231:224], a[247:240], a[255:248], a[263:256], a[271:264], a[279:272], a[287:280], a[303:296], a[311:304], a[319:312], a[327:320], a[335:328], a[343:336], a[359:352], a[367:360], a[375:368], a[383:376], a[391:384]}, w1);
matdet6 md2({a[63:56], a[71:64], a[87:80], a[95:88], a[103:96], a[111:104], a[119:112], a[127:120], a[143:136], a[151:144], a[159:152], a[167:160], a[175:168], a[183:176], a[199:192], a[207:200], a[215:208], a[223:216], a[231:224], a[239:232], a[255:248], a[263:256], a[271:264], a[279:272], a[287:280], a[295:288], a[311:304], a[319:312], a[327:320], a[335:328], a[343:336], a[351:344], a[367:360], a[375:368], a[383:376], a[391:384]}, w2);
matdet6 md3({a[63:56], a[71:64], a[79:72], a[95:88], a[103:96], a[111:104], a[119:112], a[127:120], a[135:128], a[151:144], a[159:152], a[167:160], a[175:168], a[183:176], a[191:184], a[207:200], a[215:208], a[223:216], a[231:224], a[239:232], a[247:240], a[263:256], a[271:264], a[279:272], a[287:280], a[295:288], a[303:296], a[319:312], a[327:320], a[335:328], a[343:336], a[351:344], a[359:352], a[375:368], a[383:376], a[391:384]}, w3);
matdet6 md4({a[63:56], a[71:64], a[79:72], a[87:80], a[103:96], a[111:104], a[119:112], a[127:120], a[135:128], a[143:136], a[159:152], a[167:160], a[175:168], a[183:176], a[191:184], a[199:192], a[215:208], a[223:216], a[231:224], a[239:232], a[247:240], a[255:248], a[271:264], a[279:272], a[287:280], a[295:288], a[303:296], a[311:304], a[327:320], a[335:328], a[343:336], a[351:344], a[359:352], a[367:360], a[383:376], a[391:384]}, w4);
matdet6 md5({a[63:56], a[71:64], a[79:72], a[87:80], a[95:88], a[111:104], a[119:112], a[127:120], a[135:128], a[143:136], a[151:144], a[167:160], a[175:168], a[183:176], a[191:184], a[199:192], a[207:200], a[223:216], a[231:224], a[239:232], a[247:240], a[255:248], a[263:256], a[279:272], a[287:280], a[295:288], a[303:296], a[311:304], a[319:312], a[335:328], a[343:336], a[351:344], a[359:352], a[367:360], a[375:368], a[391:384]}, w5);
matdet6 md6({a[63:56], a[71:64], a[79:72], a[87:80], a[95:88], a[103:96], a[119:112], a[127:120], a[135:128], a[143:136], a[151:144], a[159:152], a[175:168], a[183:176], a[191:184], a[199:192], a[207:200], a[215:208], a[231:224], a[239:232], a[247:240], a[255:248], a[263:256], a[271:264], a[287:280], a[295:288], a[303:296], a[311:304], a[319:312], a[327:320], a[343:336], a[351:344], a[359:352], a[367:360], a[375:368], a[383:376]}, w6);
mul m0(a[7:0], w0, w7);
mul m1(a[15:8], w1, w8);
mul m2(a[23:16], w2, w9);
mul m3(a[31:24], w3, w10);
mul m4(a[39:32], w4, w11);
mul m5(a[47:40], w5, w12);
mul m6(a[55:48], w6, w13);
sub op0(w7, w8, w14);
add op1(w14, w9, w15);
sub op2(w15, w10, w16);
add op3(w16, w11, w17);
sub op4(w17, w12, w18);
add op5(w18, w13, det);
endmodule
